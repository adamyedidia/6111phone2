library verilog;
use verilog.vl_types.all;
entity randomnessExtractor_tb is
end randomnessExtractor_tb;
