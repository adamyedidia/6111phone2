library verilog;
use verilog.vl_types.all;
entity testSerial is
end testSerial;
