library verilog;
use verilog.vl_types.all;
entity receiveBit_tb is
end receiveBit_tb;
